module Question_ROM (
    input clk,
    input [13:0] address, // ??????? pixel ?????????????? (???????? x, y)
    output reg [11:0] pixel_data // ?? RGB 12-bit (4??? 4????? 4???????)
);
    // ???????????????: ?????? IP Core Block Memory Generator
    // ???????????? .coe ??????????????????
    // ????????????????? "?????" ????????????????????????????? logic ???????????
    
    // ?????: address ??????????????????? (256) ???????????
    // ???????? address ??????? pattern ?????
    
    always @(posedge clk) begin
        // --- ??????????????????????????????????? IP Core instance ---
        // ????????: ??? address ?????????????????? 1 ????????, ????? 2 ??????? ???
        // ????? test ??? id ?????????????????????????
        pixel_data <= (address[13:10] * 12'h111) + 12'h333; 
    end
endmodule