`timescale 1ns / 1ps

module Position_Counter(
    input clk_100mhz,
    input reset,
    
    // ????????????? Move Logic (???? Pulse ?????)
    input move_left,
    input move_right,
    
    // Output ????? VGA
    output reg [9:0] rope_pos_x
    );

    // --- Config Parameters ---
    localparam CENTER_X  = 10'd320; // ????????????? (640 / 2)
    localparam STEP_SIZE = 10'd40;  // ??????????????????? (40 pixels)
    localparam MAX_WIDTH = 10'd640; // ???????????

    always @(posedge clk_100mhz) begin
        if (reset) begin
            rope_pos_x <= CENTER_X; // ??????????????????????
        end 
        else begin
            // ???????????????? (Move Left)
            if (move_left) begin
                if (rope_pos_x > STEP_SIZE) 
                    rope_pos_x <= rope_pos_x - STEP_SIZE;
                else 
                    rope_pos_x <= 0; // ??????????? (Underflow protection)
            end
            // ??????????????? (Move Right)
            else if (move_right) begin
                if (rope_pos_x < (MAX_WIDTH - STEP_SIZE)) 
                    rope_pos_x <= rope_pos_x + STEP_SIZE;
                else 
                    rope_pos_x <= MAX_WIDTH; // ???????????? (Overflow protection)
            end
        end
    end

endmodule